@00000000
13054006 9305800C 13064001 13064001
13064001 B300B500 130A1000 13014006
63040000 1301B007 9300401F 130A2000
6F000000
